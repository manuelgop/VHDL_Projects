--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   08:20:48 09/30/2013
-- Design Name:   
-- Module Name:   D:/Projects_SisDigAva/P16_Counters/Counter_vtb.vhd
-- Project Name:  P16_Counters
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Counters
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY Counter_vtb IS
END Counter_vtb;
 
ARCHITECTURE behavior OF Counter_vtb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Counters
    PORT(
         Rst : IN  std_logic;
         Clk : IN  std_logic;
         Count : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal Rst : std_logic := '0';
   signal Clk : std_logic := '0';

 	--Outputs
   signal Count : std_logic_vector(3 downto 0);

   -- Clock period definitions
   constant Clk_period : time := 100 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Counters PORT MAP (
          Rst => Rst,
          Clk => Clk,
          Count => Count
        );

   -- Clock process definitions
   Clk_process :process
   begin
		Clk <= '0';
		wait for Clk_period/2;
		Clk <= '1';
		wait for Clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      -- wait for Clk_period*10;

      -- insert stimulus here 
		Rst <= '1';
		wait for Clk_period*5;
		
		Rst <= '0';
		wait for Clk_period*20;

      wait;
   end process;

END;
