----------------------------------------------------------------------------------
-- Company:   ITESM
-- Engineer:  RickWare
-- 
-- Create Date:    17:04:15 10/09/2013 
-- Design Name: Structural Clock
-- Module Name:    Clock - Behavioral 
-- Project Name: Structural Clock
-- Target Devices: Spartan 6 (Nexys 3(
-- Tool versions: ISE WebPack v14.6
-- Description:  Using Structural (Hierarchical) VHDL
--               define a military format clock that
--               counts from 00:00:00 to 23:59:59
-- Dependencies: None
--
-- Revision: v2.0 (According to the provided schematic)
-- Revision 0.01 - File Created
-- Additional Comments: Highly effective way of using VHDL 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Clock is
    Port ( HorEn     : in   STD_LOGIC;
           DecEnt    : in   STD_LOGIC_VECTOR (3 downto 0);
           MinEn     : in   STD_LOGIC;
           UniEnt    : in   STD_LOGIC_VECTOR (3 downto 0);
           Rst       : in   STD_LOGIC;
           Clk100MHz : in   STD_LOGIC;
           Seg       : out  STD_LOGIC_VECTOR (7 downto 0);
           Disp      : out  STD_LOGIC_VECTOR (3 downto 0);
           SegOut    : out  STD_LOGIC_VECTOR (7 downto 0));
end Clock;

architecture Behavioral of Clock is
  -- Components are declared next
  
  -- A 1Hz timebase signal used for seconds will be
  -- obtained from the Nexys 3 100 MHz board signal
  -- A proper way of dividing frequency will be used.
  component Clk1Hz
  port (
    Rst    : in  STD_LOGIC;
    Clk    : in  STD_LOGIC;
	 ClkOut : out STD_LOGIC);
  end component;
  
  -- 4-bit BCD (Decimal counter) counting from 0 to 9
  -- The counter will have the following attributes:
  --   1) Parallel Synchronous Load when '1'
  --   2) Enable signal that freezes count when '0'
  --   3) Asynchronous reset (Rst) when '1'
  --   4) Terminal Count Output (TCO) which will take the
  --      value of '1' when the highest count has been
  --      reached
  component Cont0a9
  port (
    Load   : in  STD_LOGIC;
	 Enable : in  STD_LOGIC;
	 Rst    : in  STD_LOGIC;
	 Clk    : in  STD_LOGIC;
	 Valor  : in  STD_LOGIC_VECTOR(3 downto 0);
	 TCO    : out STD_LOGIC;
	 Cuenta : out STD_LOGIC_VECTOR(3 downto 0));
  end component;
  
  -- Counter which will count from 0 to 5
  -- The counter will have the following attributes:
  --   1) Parallel Synchronous Load when '1'
  --   2) Enable signal that freezes count when '0'
  --   3) Asynchronous reset (Rst) when '1'
  --   4) Terminal Count Output (TCO) which will take the
  --      value of '1' when the highest count has been
  --      reached
  --  Note that the size of the counter is 4-bits even if
  --  only 3-bits are needed for counting from 0 to 5. It
  --  is designed in this way to mantain consistency
  component Cont0a5
  port (
    Load   : in  STD_LOGIC;
	 Enable : in  STD_LOGIC;
	 Rst    : in  STD_LOGIC;
	 Clk    : in  STD_LOGIC;
	 Valor  : in  STD_LOGIC_VECTOR(3 downto 0);
	 TCO    : out STD_LOGIC;
	 Cuenta : out STD_LOGIC_VECTOR(3 downto 0));
  end component;
  
  -- Counter that count from 00 to 23 (Hour counter)
  -- The counter will have the following attributes:
  --   1) Parallel Synchronous Load when '1'
  --   2) Enable signal that freezes count when '0'
  --   3) Asynchronous reset (Rst) when '1'
  component Cont0a23
  port (
    Load     : in  STD_LOGIC;
	 Enable   : in  STD_LOGIC;
	 Rst      : in  STD_LOGIC;
	 Clk      : in  STD_LOGIC;
	 ValorDec : in  STD_LOGIC_VECTOR(3 downto 0);
	 ValorUni : in  STD_LOGIC_VECTOR(3 downto 0);
	 Cuenta   : out STD_LOGIC_VECTOR(7 downto 0));
  end component;
  
  -- A 200Hz timebase signal used for demultiplexing
  -- the 7-segment displays  will be
  -- obtained from the Nexys 3 100 MHz board signal
  -- A proper way of dividing frequency will be used.
  component RefreshDisplay
  port (
    Rst    : in  STD_LOGIC;
    Clk    : in  STD_LOGIC;
	 ClkOut : out STD_LOGIC);
  end component;
  
  -- 2-bit binary counter thar will we used to select both
  -- the display's Anode and to output the proper counter 
  component Cont0a3
  port (
    Enable  : in  STD_LOGIC;
	 Rst     : in  STD_LOGIC;
	 Clk     : in  STD_LOGIC;
	 Cuenta  : out STD_LOGIC_VECTOR(1 downto 0));
  end component;
  
  -- According to the count generated by component
  -- Cont0a3 the clock counter value will be sent to
  -- the 7-segment display after being decoded
  component Mux4to1
  port (
    DecHor  : in  STD_LOGIC_VECTOR(3 downto 0);
	 UniHor  : in  STD_LOGIC_VECTOR(3 downto 0);
	 DecMin  : in  STD_LOGIC_VECTOR(3 downto 0);
	 UniMin  : in  STD_LOGIC_VECTOR(3 downto 0);
	 Sel     : in  STD_LOGIC_VECTOR(1 downto 0);
	 Tiempo  : out STD_LOGIC_VECTOR(3 downto 0));
  end component;
  
  -- According to the count generated by component
  -- Cont0a3 the clock counter value will be selecting
  -- the Anode of the 7-segment display
  component SelAnodo
  port (
    Sel     : in  STD_LOGIC_VECTOR(1 downto 0);
	 Anodo   : out STD_LOGIC_VECTOR(3 downto 0));
  end component;
  
  -- BCD (or Binary) to 7-Segment decoder
  component DecBCD7Seg
  port (
    BCD     : in  STD_LOGIC_VECTOR(3 downto 0);
	 Seg     : out STD_LOGIC_VECTOR(7 downto 0));
  end component;
  
  -- Embedded signal
  -- 1-bit embedded signals
  signal EnHoras_int    : STD_LOGIC;
  signal EnDecMin_int   : STD_LOGIC;
  signal EnUniMin_int   : STD_LOGIC;
  signal EnSeg_int      : STD_LOGIC;
  signal EnDecSeg_int   : STD_LOGIC;
  signal Clk1Hz_int     : STD_LOGIC;
  signal TCODecMin_int  : STD_LOGIC;
  signal TCOUniMin_int  : STD_LOGIC;
  signal TCODecSeg_int  : STD_LOGIC;
  signal TCOUniSeg_int  : STD_LOGIC;
  signal ClkRefresh_int : STD_LOGIC;
  
  -- 2-bit embedded signals
  signal Sel_int        : STD_LOGIC_VECTOR(1 downto 0);
  
  -- 4-bit embedded signals
  signal DecMin_int     : STD_LOGIC_VECTOR(3 downto 0);
  signal UniMin_int     : STD_LOGIC_VECTOR(3 downto 0);
  signal Tiempo_int     : STD_LOGIC_VECTOR(3 downto 0);
  
  -- 8-bit embedded signals
  signal Hor_int        : STD_LOGIC_VECTOR(7 downto 0);
  
begin
  -- Wire (Instantiate) the components
  U1 : Clk1Hz
  port map (
    Rst    => Rst,
	 Clk    => Clk100MHz,
    ClkOut => Clk1Hz_int);
	 
  U2 : Cont0a9
  port map (
    Load   => EnSeg_int,
	 Enable => Clk1Hz_int,
	 Rst    => Rst,
	 Clk    => Clk100MHz,
	 Valor  => (others => '0'),
	 TCO    => TCOUniSeg_int,
	 Cuenta => SegOut(3 downto 0));
	 
  U3 : Cont0a5
  port map (
    Load   => EnSeg_int,
	 Enable => EnDecSeg_int,
	 Rst    => Rst,
	 Clk    => Clk100MHz,
	 Valor  => (others => '0'),
	 TCO    => TCODecSeg_int,
	 Cuenta => SegOut(7 downto 4));
	 
  U4 : Cont0a9
  port map (
    Load   => MinEn,
	 Enable => EnUniMin_int,
	 Rst    => Rst,
	 Clk    => Clk100MHz,
	 Valor  => UniEnt,
	 TCO    => TCOUniMin_int,
	 Cuenta => UniMin_int);
	 
  U5 : Cont0a5
  port map (
    Load   => MinEn,
	 Enable => EnDecMin_int,
	 Rst    => Rst,
	 Clk    => Clk100MHz,
	 Valor  => DecEnt,
	 TCO    => TCODecMin_int,
	 Cuenta => DecMin_int);
	 
  U6 : Cont0a23
  port map (
    Load      => HorEn,
	 Enable    => EnHoras_int,
	 Rst       => Rst,
	 Clk       => Clk100MHz,
	 ValorDec  => DecEnt,
	 ValorUni  => UniEnt,
	 Cuenta    => Hor_int);
	 
  U7 : RefreshDisplay
  port map (
    Rst       => Rst,
	 Clk       => Clk100MHz,
	 ClkOut    => ClkRefresh_int);
	 
  U8 : Cont0a3
  port map (
    Enable    => ClkRefresh_int,
	 Rst       => Rst,
	 Clk       => Clk100MHz,
	 Cuenta    => Sel_int);
	 
  U9: Mux4to1
  port map (
    DecHor    => Hor_int (7 downto 4),
	 UniHor    => Hor_int (3 downto 0),
	 DecMin    => DecMin_int,
	 UniMin    => UniMin_int,
	 Sel       => Sel_int,
	 Tiempo    => Tiempo_int);
	 
  U10 : SelAnodo
  port map (
    Sel       => Sel_int,
	 Anodo     => Disp);

  U11 : DecBCD7Seg
  port map (
    BCD       => Tiempo_int,
	 Seg       => Seg);
	 
  -- Gates instantiation
  EnHoras_int  <= EnDecMin_int  and TCODecMin_int and Clk1Hz_int;
  EnDecMin_int <= EnUniMin_int  and TCOUniMin_int and Clk1Hz_int;
  EnUniMin_int <= TCOUniSeg_int and TCODecSeg_int and Clk1Hz_int;
  EnSeg_int    <= HorEn         or  MinEn;
  EnDecSeg_int <= TCOUniSeg_int and                   Clk1Hz_int;

end Behavioral;









