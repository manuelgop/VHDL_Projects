----------------------------------------------------------------------------------
-- Company: ITESM
-- Engineer: Manuel Gopar
-- 
-- Create Date:    17:04:39 10/09/2013 
-- Design Name: 	 Structural Clock
-- Module Name:    Clock - Behavioral 
-- Project Name: 	 Structural Clock
-- Target Devices: Basys2
-- Tool versions:  ISE webPack 14.6v
-- Description: 	 Using Structural(Hierarchical) VHDL
					--	 Define a military format clock that
					--	 Counts
--
-- Dependencies: 
--
-- Revision:  V2.0 (According to the provided schematic)
-- Revision 0.01 - File Created
-- Additional Comments: highly effective way using VHDL
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity Clock is
    Port ( HorEn :     in  STD_LOGIC;
           DecEnt :    in  STD_LOGIC_VECTOR (3 downto 0);
           MinEn :     in  STD_LOGIC;
           UniEnt :    in  STD_LOGIC_VECTOR (3 downto 0);
           Rst :       in  STD_LOGIC;
           Clk100MHz : in  STD_LOGIC;
           Seg :       out  STD_LOGIC_VECTOR (0 to 6);
           Disp :      out  STD_LOGIC_VECTOR (3 downto 0);
           SegOut :    out  STD_LOGIC_VECTOR (7 downto 0));
end Clock;

architecture Behavioral of Clock is
--Components are declare next


--A 1Hz timebase signal used for seconds will be obtained from the basys2 100 MHz board signal
--A proper way of dividing frequency will be used
component Clk1Hz
	port (
   Rst    : in  STD_LOGIC;
   Clk    :	in  STD_LOGIC;
	ClkOut : out STD_LOGIC);
end component;


--4-bit bcd decimal conter, counting from 0 to 9
-- The counter will have the following attributes:
-- 1) Parallel Synchronous Load
-- 2) Enable signal that freezes count when '0'
-- 3) Asynchronous reset when '1'
-- 4) Terminal Count Output (TCO) which will take the 
-- value of '1' when the highest count has been reached
component Cont0a9
port(
	Load : in STD_LOGIC;
	Enable : in STD_LOGIC;
	Rst : in STD_LOGIC;
	Clk : in STD_LOGIC;
	Valor : in STD_LOGIC_VECTOR(3 downto 0);
	TCO : out STD_LOGIC;
	Cuenta : out  STD_LOGIC_VECTOR(3 downto 0));
end component;

--4-bit bcd decimal conter, counting from 0 to 5
-- The counter will have the following attributes:
-- 1) Parallel Synchronous Load
-- 2) Enable signal that freezes count when '0'
-- 3) Asynchronous reset when '1'
-- 4) Terminal Count Output (TCO) which will take the 
-- value of '1' when the highest count has been reached
--**Note that the size of the counter is 4-bits even if only
--** 3-bits are needed for counting from 0 to 5. It is designed in this way to mantein consistency
component Cont0a5
port(
	Load : in STD_LOGIC;
	Enable : in STD_LOGIC;
	Rst : in STD_LOGIC;
	Clk : in STD_LOGIC;
	Valor : in STD_LOGIC_VECTOR(3 downto 0);
	TCO : out STD_LOGIC;
	Cuenta : out  STD_LOGIC_VECTOR(3 downto 0));
end component;

--COUNTER THAT COUNTS FROM 00 TO 23 (HOUR COUNTER)
--4-bit bcd decimal conter, counting from 0 to 23
-- The counter will have the following attributes:
-- 1) Parallel Synchronous Load
-- 2) Enable signal that freezes count when '0'
-- 3) Asynchronous reset when '1'
component Cont0a23
port(
	Load : in STD_LOGIC;
	Enable : in STD_LOGIC;
	Rst : in STD_LOGIC;
	Clk : in STD_LOGIC;
	ValorDec : in STD_LOGIC_VECTOR(3 downto 0);
	ValorUni : in STD_LOGIC_VECTOR(3 downto 0);
	Cuenta : out  STD_LOGIC_VECTOR(7 downto 0));
end component;

--A 200Hz timebase signal used for demultiplexing the 7 segments display will be obtained from the tablet 100MHz board signal
--A proper way of dividing frequency will be used
component RefreshDisplay
	port (
   Rst    : in  STD_LOGIC;
   Clk    :	in  STD_LOGIC;
	ClkOut : out STD_LOGIC
	);
end component;

--2-bit binary counter that will be used to select both
-- the displays anode and to output the proper counter
component Cont0a3
	port (
   Enable    : in  STD_LOGIC;
   Rst    :	in  STD_LOGIC;
	Clk : in STD_LOGIC;
	Cuenta : out STD_LOGIC_VECTOR( 1 downto 0));
end component;


--According to the count generated by component 
--Count0a3 the.... 
component Mux4to1
	port (
   DecHor    : in  STD_LOGIC_VECTOR( 3 downto 0);
   UniHor    :	in  STD_LOGIC_VECTOR( 3 downto 0);
	DecMin :	in  STD_LOGIC_VECTOR( 3 downto 0);
	UniMin :	in  STD_LOGIC_VECTOR( 3 downto 0);
	Sel :	in  STD_LOGIC_VECTOR( 1 downto 0);
	Tiempo :	out  STD_LOGIC_VECTOR( 3 downto 0));
end component;


--According to the count generated by componene 
--Cont0a3 the clock counter value will be selecting 
-- the anode of the 7-segment display
component SelAnodo 
	port(
	Sel :	in  STD_LOGIC_VECTOR( 1 downto 0);
	Anodo :	out  STD_LOGIC_VECTOR( 3 downto 0));
end component;


--BCD(OR BINARY) to 7-segment decoder
component DecBCD7Seg 
	port(
	BCD :	in  STD_LOGIC_VECTOR( 3 downto 0);
	Seg :	out  STD_LOGIC_VECTOR( 0 to 6));
end component;


--EMBEDDED SIGNALS
--1-bit embedded signals
signal EnHoras_int : STD_LOGIC;
signal EnDecMin_int : STD_LOGIC;
signal EnUniMin_int : STD_LOGIC;
signal EnSeg_int : STD_LOGIC;
signal EnDecSeg_int : STD_LOGIC;
signal Clk1Hz_int : STD_LOGIC;
signal TCODecMin_int : STD_LOGIC;
signal TCOUniMin_int : STD_LOGIC;
signal TCODecSeg_int : STD_LOGIC;
signal TCOUniSig_int : STD_LOGIC;
signal ClkRefresh_int : STD_LOGIC;


--2-bits embedded signals
signal Sel_int : STD_LOGIC_VECTOR (1 downto 0);
--4-bits embedded signals
signal DecMin_int : STD_LOGIC_VECTOR (3 downto 0);
signal UniMin_int : STD_LOGIC_VECTOR (3 downto 0);
signal Tiempo_int : STD_LOGIC_VECTOR (3 downto 0);

--8-bits embedded sinal
signal Hor_int : STD_LOGIC_VECTOR (7 downto 0);

begin
--WIRE(Instantiate) the components

U1 : Clk1Hz
port map (
   Rst => Rst,
	Clk => Clk100Mhz,
	ClkOut => Clk1Hz_int);

U2 : Cont0a9
port map (
	Load => EnSeg_int,
	Enable => Clk1Hz_int,
	Rst => Rst,
	Clk => Clk100MHz,
	Valor => (others => '0'),
	TCO => TCOUniSig_int,
	Cuenta => SegOut (3 downto 0));
	
U3 : Cont0a5
port map (
	Load => EnSeg_int,
	Enable => EnDecSeg_int,
	Rst => Rst,
	Clk => Clk100MHz,
	Valor => (others => '0'),
	TCO => TCODecSeg_int,
	Cuenta => SegOut (7 downto 4));

U4 : Cont0a9
port map (
	Load => MinEn,
	Enable => EnUniMin_int,
	Rst => Rst,
	Clk => Clk100MHz,
	Valor => UniEnt,
	TCO => TCOUniMin_int,
	Cuenta => UniMin_int);
	
U5 : Cont0a5
port map (
	Load => MinEn,
	Enable => EnDecMin_int,
	Rst => Rst,
	Clk => Clk100MHz,
	Valor => DecEnt,
	TCO => TCODecMin_int,
	Cuenta => DecMin_int);


U6 : Cont0a23
port map (
	Load => HorEn,
	Enable => EnHoras_int,
	Rst => Rst,
	Clk => Clk100MHz,
	ValorDec => DecEnt,
	ValorUni => UniEnt,
	Cuenta => Hor_int);


U7 : RefreshDisplay
port map (
	Rst => Rst,
	Clk => Clk100MHz,
	ClkOut => ClkRefresh_int);
	
	
U8 : Cont0a3
port map (
	Enable => ClkRefresh_int,
	Rst => Rst,
	Clk => Clk100MHz,
	Cuenta => Sel_int);
	
U9 : Mux4to1
port map (
	DecHor => Hor_int (7 downto 4),
	UniHor => Hor_int (3 downto 0),
	DecMin => DecMin_int,
	UniMin => UniMin_int,
	Sel => Sel_int,
	Tiempo => Tiempo_int);
	
U10 : SelAnodo
port map(
	Sel => Sel_int,
	Anodo => Disp);
	
U11 : DecBCD7seg
port map(
	BCD => Tiempo_int,
	Seg => Seg);
	
	
	
	
	--GATES INSTANTIATION
	EnHoras_int <= EnDecMin_int and TCODecMin_int and Clk1Hz_int;
	EnDecMin_int <= EnUniMin_int and TCOUniMin_int and Clk1Hz_int;
	EnUnimin_int <= TCOUniSig_int and TCODecSeg_int and Clk1Hz_int;
	EnSeg_int <= HorEn or MinEn;
	EnDecSeg_int <= TCOUniSig_int and Clk1Hz_int;--sig seg
	
end Behavioral;
